`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Universidade Federal do Cear�
// Engineer: Lucas Esteves Rocha
// 
// Create Date: 01.08.2018 21:57:42
// Module Name: HelloWorld
// Project Name: Verilog Course
// Revision 0.01 - File Created
// 
//////////////////////////////////////////////////////////////////////////////////


module HelloWorld;
    initial begin
    $display("Hello World");
    end
    
endmodule
